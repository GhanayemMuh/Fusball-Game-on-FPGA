// (c) Technion IIT, Department of Electrical Engineering 2021 
// updated Rana Shbat May 2022


module	LevelsBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic	[1:0] level_two,
					
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout //rgb value from the bitmap  
 );

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 4;  // 2^4 = 16 
localparam  int OBJECT_NUMBER_OF_X_BITS = 6;  // 2^6 = 64 

localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


// note: sometimes, if you get a bad picture useing the MATLAB bitmap generator code
// you have to switch the X and Y sizes 

logic [0:2][0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] Levels = {{
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'h92, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'h92, 8'h92, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'h92, 8'hFF, 8'hDB, 8'h92, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h92, 8'hDB, 8'hFF, 8'hDB, 8'h92, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'h92, 8'hDB, 8'hFF },
{8'h6E, 8'h96, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h96, 8'h96, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFB, 8'h72, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h96, 8'h72, 8'hFF, 8'h96, 8'h72, 8'h96, 8'h96, 8'h72, 8'h72, 8'h72, 8'h72, 8'h96, 8'hFF, 8'hDA, 8'h72, 8'h92, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'h72, 8'h96, 8'h72, 8'hB6, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'h96, 8'h92, 8'h92, 8'h92, 8'hB6, 8'hFF, 8'h96, 8'h96, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h96, 8'h96, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h92, 8'h96, 8'h92, 8'h92, 8'h92, 8'hDA, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h72, 8'h96, 8'h97, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h6E, 8'h96, 8'h92, 8'h97, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hDB, 8'hDB, 8'hFF, 8'h96, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h4E, 8'hDB, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h96, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'h72, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h92, 8'h92, 8'h92, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h96, 8'hB6, 8'hDA, 8'h72, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h92, 8'h92, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'h72, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h96, 8'h92, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h72, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hFF },
{8'h72, 8'h97, 8'h96, 8'h92, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hDB, 8'h72, 8'h97, 8'h96, 8'h92, 8'h72, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'h97, 8'h97, 8'h72, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h92, 8'h92, 8'h72, 8'h92, 8'h72, 8'hB6, 8'hFF, 8'hDA, 8'h72, 8'h97, 8'h96, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hDB, 8'h72, 8'h96, 8'h72, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h92, 8'h96, 8'h97, 8'h97, 8'h92, 8'h72 },
{8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hB6, 8'hDB, 8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h72, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h92, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDA, 8'hDB, 8'h6E, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'hB6, 8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72 },
{8'hDB, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDA, 8'hFF, 8'hFF, 8'hDB, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDA, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hBA, 8'hBA, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDA, 8'hDF, 8'hFF, 8'hFF, 8'hDB, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDA, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB }
},
{
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h72, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hFF, 8'h92, 8'h72, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hB6, 8'h72, 8'h92, 8'h92, 8'h92, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'h72, 8'h72, 8'h72, 8'h92, 8'hB6, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h6E, 8'hDB, 8'h92, 8'h96, 8'h72, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h96, 8'h92, 8'hFF, 8'h72, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h72, 8'h6E, 8'hFF, 8'hFF, 8'h72, 8'h96, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h96, 8'h97, 8'h97, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h96, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hFF, 8'hB6, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'h92, 8'h97, 8'h96, 8'h92, 8'h92, 8'h92, 8'h92, 8'h96, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'h92, 8'h96, 8'h97, 8'h96, 8'h92, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'hDB, 8'hFF, 8'hFF, 8'h96, 8'h97, 8'h97, 8'h72, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h97, 8'h72, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h92, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hB6, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h96, 8'h92, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h96, 8'hB6, 8'hDB, 8'hDA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h92, 8'hB6, 8'hDB, 8'h72, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDA, 8'hDA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h96, 8'h96, 8'hB6, 8'h92, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h97, 8'h72, 8'hDA, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h92, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDA, 8'hDB, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h96, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h96, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'h96, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h72, 8'h97, 8'h97, 8'h72, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hBA, 8'hDB, 8'h72, 8'h96, 8'h72, 8'hFF, 8'hB6, 8'h72, 8'h97, 8'h97, 8'h96, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hB6 },
{8'hDB, 8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'h92, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'hFF, 8'hB6, 8'h6E, 8'h92, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hB6 },
{8'hFF, 8'hDA, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF }
},
{
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h72, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h72, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hFF, 8'h92, 8'h72, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hB6, 8'h72, 8'h92, 8'h92, 8'h92, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'h72, 8'h72, 8'h72, 8'h92, 8'hB6, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h6E, 8'hDB, 8'h92, 8'h96, 8'h72, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h96, 8'h92, 8'hFF, 8'h72, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h72, 8'h6E, 8'hFF, 8'hFF, 8'h72, 8'h96, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h96, 8'h97, 8'h97, 8'h96, 8'h72, 8'hBA, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h96, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'hFF, 8'hB6, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h92, 8'hB6, 8'hFF, 8'h92, 8'h97, 8'h96, 8'h92, 8'h92, 8'h92, 8'h92, 8'h96, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'h92, 8'h96, 8'h97, 8'h96, 8'h92, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'hDB, 8'hFF, 8'hFF, 8'h96, 8'h97, 8'h97, 8'h72, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h97, 8'h72, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hDA, 8'h72, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h97, 8'h92, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h96, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h96, 8'hB6, 8'hDB, 8'hDA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h92, 8'hB6, 8'hDB, 8'h72, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDA, 8'hDA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h97, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h72, 8'h96, 8'h96, 8'hB6, 8'h92, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h92, 8'h92, 8'h96, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hDB, 8'hDB, 8'hFF, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDA, 8'hDB, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hB6, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h92, 8'hDA, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'h72, 8'h6E, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF },
{8'hDB, 8'h72, 8'h97, 8'h96, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'h96, 8'h97, 8'h97, 8'h92, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h72, 8'h97, 8'h97, 8'h72, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'h72, 8'h97, 8'h97, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hBA, 8'hDB, 8'h72, 8'h96, 8'h72, 8'hFF, 8'hB6, 8'hB6, 8'hB6, 8'h96, 8'h96, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hFF },
{8'hDB, 8'h6E, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'h92, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hFF, 8'hFF, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h6E, 8'hB6, 8'hDB, 8'h6E, 8'h72, 8'h92, 8'hFF, 8'hB6, 8'hB6, 8'hB6, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'h72, 8'hFF },
{8'hFF, 8'hDA, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hDB, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hFF }
}
};

// pipeline (ff) to get the pixel color from the array 	 
//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'hFF;
	end
	else begin

		if (InsideRectangle == 1'b1 )begin  // inside an external bracket 
				RGBout <= Levels[level_two-1][offsetY][offsetX];		
		end		
//			RGBout <=  {HitEdgeCode, 4'b0000 } ;  //get RGB from the colors table, option  for debug 
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule
