// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	TeamMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					//input logic random_hart,
					input logic key6IsPressed,
					input logic key4IsPressed,
					input logic maxRotate4,
					input logic maxRotate6,


					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h09 ;// RGB value in the bitmap representing a transparent pixel
int playersPos = 0;

 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 


logic [0:15] [0:15]  MazeBiMapMask= 
{16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000100000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000010000,
16'b	0000000100000001,
16'b	0000000000000000,
16'b	0000000000010000,
16'b	0000000000000000,
16'b	0000000100000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000};
 
 
 logic [0:4] [0:31] [0:31] [7:0]  object_colors  = {

   {{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h51,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h91,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h53,8'h53,8'h5a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h5b,8'h53,8'h52,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h11,8'h52,8'h52,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h52,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h11,8'h12,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h53,8'h5b,8'h5a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h5a,8'h9a,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd1,8'hd1,8'hd1,8'h91,8'h91,8'h91,8'h91,8'hd1,8'hd1,8'hd1,8'h91,8'h91,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd1,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'h91,8'h91,8'h91,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h91,8'hda,8'hda,8'h91,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'h91,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'h91,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hd9,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'h91,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'h49,8'h49,8'h89,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'h89,8'h49,8'h49,8'h49,8'h49,8'h89,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'hd2,8'hda,8'hda,8'hda,8'hd2,8'h40,8'hda,8'hda,8'hda,8'h92,8'h49,8'hda,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hc9,8'h89,8'h49,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h49,8'hc0,8'hd2,8'hd2,8'hd2,8'hd1,8'hd2,8'hda,8'hda,8'hd2,8'hd2,8'hda,8'hd2,8'hd1,8'hda,8'hda,8'hd2,8'hd2,8'hd2,8'hc0,8'hc0,8'hc0,8'h80,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h48,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hda,8'h91,8'h91,8'h91,8'h91,8'h91,8'hd1,8'h91,8'hda,8'hda,8'hda,8'hd1,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc1,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h48,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc1,8'h09,8'h09,8'h09},
	{8'h09,8'h91,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h09,8'h09,8'h09},
	{8'h09,8'hda,8'hd9,8'hd9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd9,8'hd9,8'hd9,8'hc0,8'h09,8'h09},
	{8'h09,8'h09,8'hd8,8'hd9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd9,8'hd8,8'hd9,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hd1,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'hc0,8'h80,8'h89,8'h09,8'hc0,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h49,8'h09,8'h09,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h52,8'h09,8'h09,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h9b,8'hdb,8'h09,8'h9b,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h9b,8'hdb,8'hdb,8'hdb,8'h9b,8'h9b,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'h9b,8'hdb,8'h9b,8'hdb,8'hdb,8'h9b,8'hdb,8'h09,8'h09,8'h09}}
	,
	


	{{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h11,8'h12,8'h52,8'h09,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h5b,8'h12,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd9,8'h53,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'h5a,8'h9a,8'h9a,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'hd9,8'hd9,8'h5a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hda,8'h9a,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h11,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'hd9,8'hd8,8'hd9,8'hd9,8'hd1,8'hd1,8'hd1,8'hd1,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd9,8'hd9,8'hd1,8'hd1,8'h91,8'hda,8'hda,8'hda,8'hda,8'h92,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h53,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd1,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h49,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h53,8'h5b,8'h5b,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd1,8'hd1,8'hda,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h5b,8'h5b,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h09,8'h49,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h53,8'h5b,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd1,8'hd1,8'hda,8'h89,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'h49,8'h91,8'h09,8'h09,8'h09},
	{8'h09,8'h53,8'h5b,8'h5b,8'hda,8'hd9,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'h49,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hd0,8'hd9,8'h09,8'h09},
	{8'h09,8'h12,8'h5b,8'h9a,8'hd9,8'hd9,8'hd1,8'h91,8'hda,8'hda,8'hda,8'hda,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hd9,8'hd9,8'hd9,8'hd9,8'h09},
	{8'h09,8'h5b,8'h5b,8'hd9,8'hd8,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd9,8'hda,8'h09},
	{8'h09,8'h09,8'h5a,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd8,8'hd9,8'h09},
	{8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hda,8'h91,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hda,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd9,8'hd9,8'hd9,8'h09,8'h09},
	{8'h09,8'h09,8'h11,8'hd9,8'hd1,8'hd2,8'hda,8'h00,8'h49,8'hda,8'hda,8'hda,8'hda,8'h40,8'h00,8'h00,8'hd2,8'hda,8'hda,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hc0,8'hc0,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h51,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h40,8'h00,8'hda,8'hda,8'hda,8'hd1,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h49,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'hda,8'hda,8'hda,8'h91,8'hd1,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'hd2,8'hda,8'hd1,8'hd2,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hda,8'hd1,8'hd2,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h49,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd2,8'hd2,8'hda,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h49,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc9,8'hc9,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h49,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'h49,8'h09,8'h00,8'h49,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'h80,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc9,8'hd9,8'hd9,8'hc8,8'hd1,8'h80,8'hc0,8'hc0,8'h80,8'h80,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h80,8'h80,8'h80,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h00,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h51,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09}}
	,
	
	{{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h5b,8'h12,8'h52,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h53,8'h53,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h91,8'hd9,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h5a,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'hd9,8'hd1,8'hd1,8'hd9,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'hd9,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'h91,8'hda,8'hda,8'hd2,8'hda,8'hd1,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'h91,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h92,8'hda,8'h91,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h48,8'hda,8'hda,8'h91,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h89,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'hc8,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h09},
	{8'h09,8'h09,8'hd9,8'hd9,8'hc8,8'h80,8'hc0,8'hc0,8'hc1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h48,8'h92,8'hda,8'h91,8'hd1,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h09},
	{8'h09,8'h09,8'hd9,8'hd9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'h91,8'h91,8'h00,8'h00,8'h48,8'hda,8'hda,8'hda,8'hda,8'h49,8'h00,8'hda,8'hda,8'hda,8'hd9,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h52},
	{8'h09,8'h11,8'hd9,8'hc8,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hd2,8'hda,8'hd2,8'hda,8'h00,8'h48,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hd9,8'hd8,8'h9a,8'h5b,8'h5b,8'h5b,8'h09},
	{8'h09,8'h09,8'h09,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd1,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h11},
	{8'h09,8'h09,8'h49,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hda,8'hd1,8'hd1,8'hda,8'hd2,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h12,8'h09},
	{8'h09,8'h09,8'h80,8'hc1,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hda,8'hd1,8'hd1,8'hda,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h09},
	{8'h49,8'h09,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc9,8'hda,8'hd1,8'hd1,8'hda,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'h9a,8'h5b,8'h09,8'h09},
	{8'h49,8'h00,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc9,8'hda,8'hd1,8'hda,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'h9a,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h00,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hc0,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h00,8'h80,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hda,8'hd2,8'h91,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h00,8'h80,8'hc0,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd2,8'hc9,8'hd1,8'hda,8'h91,8'h09,8'h9a,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h00,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h00,8'h09,8'h89,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h00,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h00,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd1,8'hd9,8'hc8,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h00,8'h80,8'hc0,8'hc0,8'hc0,8'hc8,8'hd9,8'hd9,8'hd9,8'hd9,8'hc8,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h00,8'h80,8'hc0,8'hc0,8'hc8,8'hd9,8'hd9,8'hd9,8'hd9,8'hc8,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h49,8'h00,8'h80,8'h81,8'hc0,8'hd9,8'hd8,8'hd9,8'hd9,8'hd1,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h00,8'h09,8'h09,8'h09,8'hd9,8'hda,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09}}
	
	,
	
	
	
	

	
	{{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h5b,8'h5b,8'h5b,8'hd9,8'hd9,8'h91,8'hda,8'h09,8'h09,8'h09,8'h09,8'h49,8'hc1,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd8,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h53,8'h53,8'h5b,8'h5b,8'hda,8'hd9,8'hd0,8'hda,8'hda,8'h91,8'h91,8'h09,8'h49,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'hd9,8'hc9,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hd2,8'hd1,8'h91,8'h89,8'hc0,8'hc0,8'hc0,8'hc0,8'hd0,8'hd9,8'hd9,8'hd0,8'hc8,8'h09,8'h92,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h12,8'h5b,8'h5b,8'h5b,8'h5b,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd9,8'hd9,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h5b,8'h5a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h5b,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h53,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h5a,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hd1,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'hd1,8'hda,8'h00,8'h00,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h09,8'h09,8'h09},
	{8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h89,8'h48,8'hd2,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09},
	{8'h48,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'h49,8'hd2,8'hd2,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h81,8'h41,8'h49,8'h09},
	{8'h09,8'h51,8'h5a,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'h49,8'hda,8'hd2,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h53,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h48,8'h49,8'hda,8'hd2,8'h91,8'hda,8'h80,8'h80,8'h80,8'h80,8'h80,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h49,8'h49,8'hda,8'hda,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h89,8'h48,8'hda,8'h91,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h52,8'h5b,8'h5b,8'h5a,8'hd9,8'hd9,8'hd1,8'hda,8'h00,8'h00,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hd1,8'hda,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h12,8'h5b,8'h5a,8'hd9,8'hd9,8'hd1,8'hda,8'hd2,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h5b,8'h9a,8'hd9,8'hd1,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h52,8'h52,8'h91,8'hd9,8'hd1,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h89,8'h40,8'h49,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h09,8'h49,8'h49,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'hda,8'hda,8'hda,8'h91,8'h09,8'h09,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hd9,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hc0,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09}}
	,
	
	{{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hda,8'h92,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd8,8'hd9,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hd9,8'hc0,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd1,8'hc0,8'hc0,8'h80,8'hc0,8'hc0,8'h09,8'h09,8'hd2,8'hda,8'hda,8'hda,8'h92,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h09,8'h09,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h01,8'h40,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h5a,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h01,8'h40,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hd1,8'hd9,8'h9a,8'h5b,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h91,8'h91,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h12,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h00,8'h00,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'h00,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h11,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'hda,8'h00,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'h80,8'h80,8'h80,8'h80,8'h80,8'hda,8'h91,8'hda,8'hda,8'h00,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'hda,8'h00,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'h51,8'h09},
	{8'h09,8'h49,8'h49,8'h81,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'h92,8'h49,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'h51},
	{8'h09,8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'h00,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hd2,8'hd2,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9},
	{8'h09,8'h09,8'h09,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h00,8'h00,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'hd9,8'hd9},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h9a,8'h91,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h5b,8'h52,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd8,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h5b,8'h11,8'h09,8'h09,8'h09},
	{8'h09,8'h00,8'h40,8'hc0,8'hc0,8'hc8,8'hd9,8'hd9,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hd1,8'hd2,8'hda,8'hda,8'hda,8'hda,8'hda,8'hd1,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hc8,8'hd1,8'hd9,8'hd9,8'hd1,8'hc0,8'hc0,8'hc0,8'hc0,8'h49,8'h91,8'hd1,8'hd1,8'hda,8'hd2,8'hd1,8'hd9,8'hd9,8'h9a,8'h5b,8'h5b,8'h5b,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hd1,8'hd9,8'hd9,8'hd9,8'hd9,8'hc0,8'hc0,8'hc0,8'h88,8'h09,8'h09,8'h91,8'h91,8'hda,8'hd1,8'hd1,8'hd9,8'h9a,8'h5b,8'h5b,8'h52,8'h52,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h9a,8'hd8,8'hd9,8'hd9,8'hd9,8'hc0,8'hc0,8'hc1,8'h09,8'h09,8'h09,8'h09,8'h51,8'hd2,8'h91,8'hd9,8'hd9,8'h5b,8'h5b,8'h5b,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'hda,8'hd9,8'hd9,8'hd9,8'hd9,8'hc0,8'hc1,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'hd9,8'hd9,8'hc0,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09}}};
 
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		playersPos <= 0;

	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		if (key6IsPressed == 1'b1) begin

			if (maxRotate6)
				playersPos <= 3;
			else
			playersPos <= 1;
		end // key6
		
		else if (key4IsPressed == 1'b1) begin
			if (maxRotate4) begin
				playersPos <= 4;
			end 
			else
				playersPos <= 2;
		end // key4
		
		else begin
			playersPos <= 0;
		end
		
		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
			(MazeBiMapMask[offsetY[8:5] ][offsetX[8:5]] == 1'b1 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[playersPos][offsetY[4:0]][offsetX[4:0]] ; 
		

	end // main else
end // ff

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

